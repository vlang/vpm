module models

pub struct Category {
pub:
	id   int
	slug string
	name string
}
