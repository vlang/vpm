module models

pub struct Category {
pub:
	id          int
	name        string
	packages int
}
