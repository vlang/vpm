module session

