module models

pub struct Tag {
pub:
	id   int
	slug string
	name string
}
