module dto

pub struct User {
pub:
	gh_id        int
	login        string
	avatar       string
	name         string
	access_token string
}
