module auth
