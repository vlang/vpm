module models

// Formatting for Postgres to_char() function
const iso8601 = 'YYYY-MM-DD"T"HH24:MI:SSOF'
