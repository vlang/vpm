module github

// !!! DO NOT USE IN YOUR PROJECT
// vpm.github implements only specific for vpm parts of api
