module models

pub struct Tag {
pub:
	id       int
	name     string
	packages int
}
