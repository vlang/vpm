module app

import web
import json

['/api/user/:login'; get]
fn (mut app App) api_user(login string) web.Result {
	user := app.services.users.get_by_login(login) or { return wrap_service_error(mut app, err) }

	return app.json(.ok, json.encode(user))
}

['/api/bans/:login'; post]
fn (mut app App) api_admin_create_user_ban(login string) web.Result {
	if !app.authorized() {
		return app.send_status(.unauthorized)
	}

	if !app.user.is_admin {
		return app.send_status(.forbidden)
	}

	user := app.services.users.get_by_login(login) or { return wrap_service_error(mut app, err) }

	app.services.users.set_blocked(user.id, true) or { return wrap_service_error(mut app, err) }

	return app.send_status(.ok)
}

['/api/bans/:login'; delete]
fn (mut app App) api_admin_delete_user_ban(login string) web.Result {
	if !app.authorized() {
		return app.send_status(.unauthorized)
	}

	if !app.user.is_admin {
		return app.send_status(.forbidden)
	}

	user := app.services.users.get_by_login(login) or { return wrap_service_error(mut app, err) }

	app.services.users.set_blocked(user.id, false) or { return wrap_service_error(mut app, err) }

	return app.send_status(.ok)
}
