module storage

pub const (
	err_not_found = error('file not found')
)
