module models

pub struct GHToken {
pub:
	user_id int
	token   string
}
