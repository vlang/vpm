module main

pub fn (mut app App) logged_in() bool {
	return false
}