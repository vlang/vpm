module log

import x.json2 as j2

struct Field {
	key string
	value j2.Any
}
