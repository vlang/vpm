module dto

pub struct User {
pub:
	gh_id           int
	gh_login        string
	gh_avatar       string
	name            string
	gh_access_token string
}
