module repository

const (
	categories_table          = 'category'
	packages_table            = 'package'
	tags_table                = 'tag'
	tokens_table              = 'token'
	users_table               = 'user'
	versions_table            = 'version'

	dependencies_table        = 'dependency'
	package_to_category_table = 'package_to_category'
	package_to_tag_table      = 'package_to_tag'
)
