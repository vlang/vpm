module models

pub struct Token {
pub:
	user_id string
	access_token string
}
