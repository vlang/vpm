module auth