module dto

pub struct User {
pub:
	gh_id    int
	gh_login string
	name string
	gh_avatar string
	gh_access_token string
}
