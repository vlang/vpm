module session
